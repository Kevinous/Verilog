

module HalfAdd(x, y, out);  
 
    input x, y;  
 
    output [1 : 0] out;  
 
    assign out = x + y;  
 
endmodule  